
module alarm_qsys (
	clk_clk,
	hex4_export,
	hex3_export,
	hex2_export,
	hex1_export,
	hex0_export,
	hex5_export,
	key_export);	

	input		clk_clk;
	output	[6:0]	hex4_export;
	output	[6:0]	hex3_export;
	output	[6:0]	hex2_export;
	output	[6:0]	hex1_export;
	output	[6:0]	hex0_export;
	output	[7:0]	hex5_export;
	input	[3:0]	key_export;
endmodule
